*AD834 Macro-model
*Function:Multiplier
*
*Revision History:
*Rev.1 Feb 2015-Initials
*Copyright 2015 by Analog Devices
*
*Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spicemodels/license
*for License Statement. Use of this model indicates your acceptance
*of the terms and provisions in the License Statement.
*
*
*Not modeled:
*	Output biasing functionality
*
*Parameters modeled include:
*   Vos, Ibias, input clipping voltage,CMRR
*   Bandwidth
*
* Node assignments
*             Y1
*             |  Y2
*             |  | -Vs
*             |  |  |  W2   
*             |  |  |  | W1  
*             |  |  |  |  | +Vs  
*             |  |  |  |  |  |  X1  
*             |  |  |  |  |  |  | X2
*             |  |  |  |  |  |  |  |   
*.SUBCKT AD834 Y1 Y2 50 W2 W1 99 X1 X2
*$
.SUBCKT AD834 Y1 Y2 VS- W2 W1 VS+ X1 X2
**********
Rx1 19 0 10000G
Rx2 5 0 10000G
Rx3 8 0 10000G
Rx4 15 0 10000G
Rx5 17 0 10000G


R18 X1 4 1 
D14 4 11 Diode
V26 11 X2 1.3 
D13 20 4 Diode
V23 X2 20 1.3
I2 X2 0 4.5e-005
I1 4 0 4.5e-005
R2 6 X2 12500
R1 4 6 12500 
E17 4 3 10 0 1
C2 9 10 3.1e-011
R4 9 10 3830 
R3 0 10 1
*
E2 9 0 6 0 1
V1 3 21 5e-005
C3 0 Xout 2.653e-016
R5 0 Xout 1000000 
G3 0 Xout 21 X2 1e-006
V13 45 VS_in- 1 
D5 45 Xout Diode
V11 VS_in+ 43 1 
D4 Xout 43 Diode
************
R25 Y1 14 1 
D7 14 29 Diode
V20 29 Y2 1.3
D6 18 14 Diode
V16 Y2 18 1.3
I5 Y2 0 4.5e-005
I4 14 0 4.5e-005
E12 14 37 28 0 1
C1 27 28 3.1e-011
R10 27 28 3830 
R9 0 28 1
E9 27 0 26 0 1
R8 26 Y2 12500 
R7 14 26 12500 
V8 37 16 5e-005 
C4 0 Yout 2.653e-016
R11 0 Yout 1000000 
G6 0 Yout 16 Y2 1e-006
V24 33 VS_in-  1 
D8 33 Yout Diode
V18 VS_in+ 30 1 
D3 Yout 30 Diode
************
E6 xy_out 0 VALUE={ V(Xout)*V(Yout) }
V31 35 VS_in- 1 
D10 35 out Diode
V30 VS_in+ 31 1 
D9 out 31 Diode
C6 0 out 3.183e-011
R34 0 out 1 
G14 0 out xy_out 19 1
R19 2 24 1000 
R17 12 48 1000 
R15 8 15 1000   
R14 5 17 1000 
E25 5 8 out 19 1
E22 0 2 17 15 1
E14 12 0 17 15 1
I10 W2 0 0.0085 
I9 W1 0 0.0085
R23 0 W2 1000000
R22 W1 0 1000000 
G8 W2 0 24 0 0.004
G7 W1 0 48 0 0.004
V35 36 VS_in- 0.5 
D15 36 W2 Diode
V34 VS_in+ 13 0.5 
D12 W2 13 Diode
V33 22 VS_in- 0.5
D11 22 W1 Diode
V29 VS_in+ 1 0.5 
D2 W1 1 Diode
*********
E3 VS_in+ mid VS+ mid 1
E4 mid VS_in- mid VS- 1
E1 mid 0 7 0 1
R13 7 VS- 10000000 
R12 VS+ 7 10000000 
.model Diode  D
.ENDS
*$
